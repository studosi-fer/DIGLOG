/* Verilog model created from schematic test2.sch -- Oct 26, 2015 01:06 */

module test2;




endmodule // test2
