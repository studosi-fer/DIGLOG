/* Verilog model created from schematic Test1.sch -- Oct 26, 2015 01:06 */

module Test1;




endmodule // Test1
