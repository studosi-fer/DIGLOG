
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library xp2;
use xp2.components.all;

--
-- Podesite generic parametar C_JMBAG!
--
-- Nije potrebno ni dozvoljeno raditi bilo kakve druge preinake u VHDL kodu!
--

entity pogodi_bistabil is
    generic (
	C_JMBAG: integer := 0012345678
    );
    port (
	btn_left, btn_center, btn_right, btn_up, btn_down: in std_logic;
	sw: in std_logic_vector(3 downto 0);
	led: out std_logic_vector(7 downto 0);
	clk_25m: in std_logic
    );
end pogodi_bistabil;

architecture x of pogodi_bistabil is
    signal d, e, s, r, j, k, t, clk: std_logic;
    signal q: std_logic_vector(7 downto 0);

    -- Ovo treba samo za debouncing signala takta (clk)
    signal clk_cnt: integer;

    -- Ovo treba samo za hash mux:
    signal addr_a, addr_b: std_logic_vector(12 downto 2);
    signal data_a, data_b: std_logic_vector(31 downto 0);
    signal pre_mask: std_logic_vector(7 downto 0);

begin
    -- clk je upravljan tipkom "btn_right" preko debouncing sklopa
    d <= btn_left;
    e <= btn_center;
    s <= btn_up;
    r <= btn_down;
    j <= btn_up;
    k <= btn_down;
    t <= btn_left;

    --
    -- "SR" bistabil
    --
    -- U tablicu upisati: SR
    --
    process(s, r)
    begin
	if s = '1' then
	    q(0) <= '1';
	elsif r = '1' then
	    q(0) <= '0';
	end if;
    end process;

    --
    -- "D" bistabil s enable ulazom (latch)
    --
    -- U tablicu upisati: D latch
    --
    process(d, e)
    begin
	if e = '1' then
	    q(1) <= d;
	end if;
    end process;

    --
    -- "D" bistabil okidan rastucim bridom takta (flip-flop)
    --
    -- U tablicu upisati: D flip-flop
    --
    process(clk)
    begin
	if rising_edge(clk) then
	    q(2) <= d;
	end if;
    end process;

    --
    -- "D" bistabil okidan rastucim bridom takta (flip-flop)
    -- i asinkronim set / reset ulazima
    --
    -- U tablicu upisati: D flip-flop, asinkroni SR
    --
    process(clk, s, r)
    begin
	if s = '1' then
	    q(3) <= '1';
	elsif r = '1' then
	    q(3) <= '0';
	elsif rising_edge(clk) then
	    q(3) <= d;
	end if;
    end process;

    --
    -- "D" bistabil okidan rastucim bridom takta (flip-flop)
    -- i sinkronim set / reset ulazima
    --
    -- U tablicu upisati: D flip-flop, sinkroni SR
    --
    process(clk)
    begin
	if rising_edge(clk) then
	    if s = '1' then
		q(4) <= '1';
	    elsif r = '1' then
		q(4) <= '0';
	    else
		q(4) <= d;
	    end if;
	end if;
    end process;

    --
    -- "D" bistabil okidan rastucim bridom takta (flip-flop) s enable ulazom
    -- i sinkronim set / reset ulazima
    --
    -- U tablicu upisati: D flip-flop s enable ulazom, sinkroni SR
    --
    process(clk)
    begin
	if rising_edge(clk) then
	    if s = '1' then
		q(5) <= '1';
	    elsif r = '1' then
		q(5) <= '0';
	    elsif e = '1' then
		q(5) <= d;
	    end if;
	end if;
    end process;

    --
    -- "T" bistabil
    --
    -- U tablicu upisati: T
    --
    process(clk)
    begin
	if rising_edge(clk) and t = '1' then
	    q(6) <= not q(6);
	end if;
    end process;

    --
    -- "JK" bistabil
    --
    -- U tablicu upisati: JK
    --
    process(j, k, clk)
    begin
	if rising_edge(clk) then
	    if j = '1' and k = '1' then
		q(7) <= not q(7);
	    elsif j = '1' then
		q(7) <= '1';
	    elsif k = '1' then
		q(7) <= '0';
	    end if;
	end if;
    end process;


    --
    -- Debouncer signala takta
    --
    -- NE DIRAJTE I NE MIJENJAJTE OVAJ DIO VHDL KODA!
    --

    process(clk_25m)
    begin
	if rising_edge(clk_25m) then
	    if btn_right /= clk then
		if clk_cnt = 250000 then -- 10 ms
		    clk <= btn_right;
		else
		    clk_cnt <= clk_cnt + 1;
		end if;
	    else
		clk_cnt <= 0;
	    end if;
	end if;
    end process;

    --
    -- Prospojnik izlaza iz bistabila na LED indikatore.
    --
    -- NE DIRAJTE I NE MIJENJAJTE OVAJ DIO VHDL KODA!
    --

    addr_a <= std_logic_vector(to_unsigned(C_JMBAG, 11));
    addr_b <= data_a(10 downto 0);

    G_iter: for i in 0 to 7 generate
    begin
	with data_b(((i * 4) + 2) downto (i * 4)) select
	pre_mask(i) <=
	    q(0) when "000",
	    q(1) when "001",
	    q(2) when "010",
	    q(3) when "011",
	    q(4) when "100",
	    q(5) when "101",
	    q(6) when "110",
	    q(7) when "111";
	led(i) <= pre_mask(i) when sw(3) = '0' or
	  to_integer(unsigned(sw(2 downto 0))) = i else '0';
    end generate;
 
	ram_8_0: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B => "NORMAL", WRITEMODE_A => "NORMAL",
		GSR => "ENABLED", RESETMODE=> "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A => "NOREG",
		DATA_WIDTH_B => 9, DATA_WIDTH_A => 9,
		INITVAL_00 => "0x192FA0B2F00B604116E511CE5052FD002711A2731FADC1308C116F414AB8096D714C0402AEA1CACA",
		INITVAL_01 => "0x018B409ECB1A276118AB1568E0B4C9180A71D8BD1C6EF184B0164AF04C960124E1808B11A370B826",
		INITVAL_02 => "0x1F486050840E6FC1BED30D09D06E3902C0D1CEBA02AB50F2291904D1D2CE12E521BE410702317E7E",
		INITVAL_03 => "0x05845184DA02A3E10A7E02C87102701FCE7102B1106F005CC31B6290909E1020C16C4A1E27201CAC",
		INITVAL_04 => "0x04E0300252114DF106920BE560E23413A250C8F20A4670F6671CA5C184490AC890A22905A841C097",
		INITVAL_05 => "0x0422115E10156BD084321FAEA0049313C47060AE0B632190A5118D40F0560B2F60E452018341A461",
		INITVAL_06 => "0x09A760D8091B00E048B70B6B909A3C072D00748E0FC7A0BC7B0482E1128F03EC61CE581B6A50FA3C",
		INITVAL_07 => "0x0EC5607016114270946F1BC8F148310DA451A205036AF0F49009C48080021802C04A3E01CF21F8C6",
		INITVAL_08 => "0x07E300F804006C6070290D8AE08C9A15038024F11EA0F0727B07E3606E930F0F310C530C6A80C6D2",
		INITVAL_09 => "0x012A71E86117E1A068051060C0DEA813AE3042CE118781BE0F0904F00848136B911CEA1D4DB06818",
		INITVAL_0a => "0x10A4A1E2E3060C01C8301BE13016C31FCE91965B0A68D08EAB0928B0261D02C4E1BC2607A181603D",
		INITVAL_0b => "0x1C6F406A500F26C1E2A618AEB1A2CF06EF4186DC164861FC42096E417CE30866D182F801AF0004E4",
		INITVAL_0c => "0x08A5602494104160D2B20EC5904E9006CBF0F8D702A02118BE0FC530627D10AAD0AE41006E415052",
		INITVAL_0d => "0x01E811521804CC2158341CA051AC9F15E39030C6174F41FAE21BC650E63F17E1806ABC13E6C0DA85",
		INITVAL_0e => "0x14A1A1A8D306E2510EC30748E11C211F6EF1146A1C68A146B111AA8068540C4510D8D90C2FE1A646",
		INITVAL_0f => "0x0301409CB50167E046071702E1F87404C8411C5F184401B28700C8B018B2018DC1A48C12EDB18239",
		INITVAL_10 => "0x006151F40106C74196900BCFA140730B2810B8EF03A3D1CE3F0302E12C1706217194FC09E4D15863",
		INITVAL_11 => "0x0702307E0F180FA0F8B11A8CD028051EAA30E0C70F2E302871092E40D0860022407C1B1948E1D62F",
		INITVAL_12 => "0x1AE28092F00B86512C450FAC503EAE00A0A0C89E050970F40F18614016F310E311AE380B83201E76",
		INITVAL_13 => "0x14C9D0CE571D87E1C09C164A41DA400B6F11EA9803894090AD0800A00AB10366A1F2C91F6E103871",
		INITVAL_14 => "0x0F80D0A4710E895018B40865B1B08F0D2301D23F120540F6461FC230B4E711A2903CBF064471B4FD",
		INITVAL_15 => "0x0021602C8B0E6A81AC16056730C63F0C23F11E8D12463018C0164960E6260748118CF91A4E71705B",
		INITVAL_16 => "0x158CB1DEB909E591D0100621417E631BC411564A0DE2B020FC0267D0C4B215A7305E5A086CE1261A",
		INITVAL_17 => "0x14C29160B20A8F211C150D4E80A2CB1CAC5128DC0DA4503AC30302607E2B1925A1406719AF819C69",
		INITVAL_18 => "0x1F04B10CC707CE30B0961621F06AEB1E6E90EAE20D8181E857108F807E79190541A6F205E030260D",
		INITVAL_19 => "0x1C2CB016500263917E521028504EE10E0171A6841145A004340060700AA1074E319A690AC3E140FB",
		INITVAL_1a => "0x1A41E058C511A9D040601F06D0CED909E4E1B0CB0E6481A82B16A791A4240A83418ED7190E41C616",
		INITVAL_1b => "0x04EA01BCB70C22707C831627B12A2E0DE760A2DB186C702A1717872102541E0D60F4B71DA2E1728B",
		INITVAL_1c => "0x1C241024281FCDB06A3113CB401CCE1F48D17C42152DE1269B1F6C8160611E243164D71E6051F27B",
		INITVAL_1d => "0x178FC168A10A89A0B613040AC07C7218AB8112210D8050E66A152BC1DA25058C71A85E04A2B19C64",
		INITVAL_1e => "0x1B232162AD18017096CE14A5E1DE6D16C32056FA0CA4116413194A50649F1FC141A42C1DEA909CF0",
		INITVAL_1f => "0x01698036FE0B4A11EA50090AE17E3C1900D1269C1C2B7180500806C140701A6F600CD61FC35170B8",
		INITVAL_20 => "0x0F89B07A70086580B282162821F2FE06E8C1EC8B160310A04E1A60119A2C194830565F00C3E18A4A",
		INITVAL_21 => "0x1B6D717CE2070C10D8CA0A62910623150AF184D91C6A41B62C008B6182FC1BC7B030981BEBD09C2B",
		INITVAL_22 => "0x1AED20908F1066B02A5F0EA9E13AA91843E1E6170AEF60C8501E0A51E25B1EA6F0BCB615EA0036CD",
		INITVAL_23 => "0x0CA9206CF512C7B12A0C15C01016FD09A4E1906306279178D118E1305828040C11B86D02E97036DE",
		INITVAL_24 => "0x0BC510EC9C1E0D01D85C196B203AAC1D2B61D2C71F01E0787D050FC0F0EA0E62B1FC7D138B404C03",
		INITVAL_25 => "0x1424617ED30281C1A6E105653114CF08AEA1C8E8050AD0E8250A09C0E0CA0FA0B14845062B00B4CF",
		INITVAL_26 => "0x1FC260D6CB11CAF00C0D0B02506C7514C620F46808E7503EE7002490E8DB056C810AC801C7316418",
		INITVAL_27 => "0x16C40092631DA731A2FB04CD90568B03EF31C697126AC15A8907A23174B012858156E101C1C094E1",
		INITVAL_28 => "0x1B0AF074D31C4A51827E186120B25A140FD02C2815A69196590F6400A84D15E2D040CD128D815234",
		INITVAL_29 => "0x0E67B1E85612C5C0A8CE1F4120122819AFE192BA068200D2650121A0B4480AC4A1E4E802ED114E59",
		INITVAL_2a => "0x07C8109AFE0EC5E0708B05C6D1C05B13E8D0B8020E6D605C451EC9C09E350527D1DEC70C4CA10498",
		INITVAL_2b => "0x17AC812CC5150691843808E1A19CAB0721703C0E1C2EA1FA351C6BF1B27E1844817C431A034138EF",
		INITVAL_2c => "0x0EA0918AC612E8504CF21720908CFB05A9D106021EC900425003C370BE6B05CEF1F4560288603045",
		INITVAL_2d => "0x16EA511CED1E85403E2E1C0F60844D0A67B0788F148780B82608EAE162AC14CD91F043024EF04A90",
		INITVAL_2e => "0x018F919E7C014F400AFD0DA07192830FA7B0129E05C410F6D0020411406D08014064140405301C68",
		INITVAL_2f => "0x004E901EE111E6309ADB1069506A351ECBF14A040DA130366219CFD19C9B0EA020BC0702646086EC",
		INITVAL_30 => "0x1C41400267028D11C839150501A2FD1C6FA018A618250060B803E7E1A4FC1CA9D1825102CAF0BCAC",
		INITVAL_31 => "0x1945600AA01D0711D6181B48E038530048B0D63C028AD06C50006AB11E9A140E5092271E24918C01",
		INITVAL_32 => "0x180180DA791B46718A0B1CA49180E8062A9060D1086300DAD21181D16EB8062381DA4F1401717CC5",
		INITVAL_33 => "0x11EEF01CA90200F03AF91367E0CA431267A07C3417A0A0B09A1047C06E640B6AF0F4950068A01658",
		INITVAL_34 => "0x04E3209CA700AA718CA50687A10C161A8FC1D00F04EDC138B51B2210FAA00B83C0B445082060B661",
		INITVAL_35 => "0x190C91AE271A8D200465082A00C0C8038600B4C5042820148D0F0B6174D419A70146571EC64192C6",
		INITVAL_36 => "0x1807A0FC8109C3E0F28D1CED00D4FB0BECB1E043072E11B01C092BE1D237094DB01E6A196C302C1F",
		INITVAL_37 => "0x0FAA806CD7070601A67B1DA8F158CE19A8A19A9A1847907C42190951F4D01DE5A1EA5106C7411E21",
		INITVAL_38 => "0x15E581C6201E2CF1E63406AAE1EC3610C9B1386D16A510E8E001ED710E4619A731E6030D8BC03643",
		INITVAL_39 => "0x0A2231C838156C81EC890CA2C01E7E17EA90487908A5009C101B8061F2360DE9D0F66B040D91EAF5",
		INITVAL_3a => "0x00C90030DB1C2820469C07ACA158D90AED6040211A8D91908C0860715A1D00C95180951269208081",
		INITVAL_3b => "0x1424F0A05616C560CEC81D2400E00516EB90387E1EA1F1384B02ED80142D17EC311A891F4A10A47C",
		INITVAL_3c => "0x128031920F1D42117E2401CEA1064D13E04168EA07AD7036A70A2A403E201A4CB09A140F2400FC5F",
		INITVAL_3d => "0x17447140EB1F4011D632150D60F0E31DA1D1921D1F2101C22714ACE0F64A17AA30400A114AE0CA6C",
		INITVAL_3e => "0x114E31368F024B8038A40A83E0622E0DA531860D04E3117EB806CA018CCA1F2811C07810A0618062",
		INITVAL_3f => "0x0DA64052EB1C42C130650E21C13E500F4530B834134D40B6141F40B18CA8084530E8F51B2AC11859"
	)
	port map (
		DIA0 => '0', DIA1 => '0', DIA2 => '0', DIA3 => '0',
		DIA4 => '0', DIA5 => '0', DIA6 => '0', DIA7 => '0',
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => data_b(0), DOA1 => data_b(1),
		DOA2 => data_b(2), DOA3 => data_b(3),
		DOA4 => data_b(4), DOA5 => data_b(5),
		DOA6 => data_b(6), DOA7 => data_b(7),
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0', ADA2 => '0', 
		ADA3 => addr_b(2), ADA4 => addr_b(3),
		ADA5 => addr_b(4), ADA6 => addr_b(5),
		ADA7 => addr_b(6), ADA8 => addr_b(7),
		ADA9 => addr_b(8), ADA10 => addr_b(9),
		ADA11 => addr_b(10), ADA12 => addr_b(11),
		ADA13 => addr_b(12),
		CEA => '1', CLKA => clk_25m, WEA => '0',
		CSA0 => '0', CSA1 => '0', CSA2 => '0', RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => data_a(0), DOB1 => data_a(1),
		DOB2 => data_a(2), DOB3 => data_a(3),
		DOB4 => data_a(4), DOB5 => data_a(5),
		DOB6 => data_a(6), DOB7 => data_a(7),
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0', ADB2 => '0', 
		ADB3 => addr_a(2), ADB4 => addr_a(3),
		ADB5 => addr_a(4), ADB6 => addr_a(5),
		ADB7 => addr_a(6), ADB8 => addr_a(7),
		ADB9 => addr_a(8), ADB10 => addr_a(9),
		ADB11 => addr_a(10), ADB12 => addr_a(11),
		ADB13 => addr_a(12),
		CEB => '1', CLKB => clk_25m, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	ram_8_1: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B => "NORMAL", WRITEMODE_A => "NORMAL",
		GSR => "ENABLED", RESETMODE => "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A=> "NOREG",
		DATA_WIDTH_B => 9, DATA_WIDTH_A => 9,
		INITVAL_00 => "0x1E0561D4421C42F1ACF20B83F17E640AC4A11894174F01E6650843D0E6E90D4431E0F505C1318059",
		INITVAL_01 => "0x04EA00D695040A01CE980029F0822D0B20401271002B80E04501E5003A350AE130C65F1F88907210",
		INITVAL_02 => "0x16AF913A360283A11C1A0E43C1A8D60F032142CD068CF06C4B1722709A571C09E01C2B0DA471D4C1",
		INITVAL_03 => "0x17C2611E340181C16C181E8D617EA3186B01CE040826D06A56052BD1EAC3046A304A071B64B07A79",
		INITVAL_04 => "0x082CD1E604092041E20E1148710C690F47B04E3D17ED912049020BE10E0B0E23A096E802CD9186C6",
		INITVAL_05 => "0x1AC6F0BC6300A761E047138450380C196B00D2D315C761A2C716A37158C10DE411AC7B12C611F278",
		INITVAL_06 => "0x140941A2BF0FCD71DEDE082860CE1F09CAC0C8A317284112C112E9D1BE9A11C75174130F4C911C9F",
		INITVAL_07 => "0x12A1B134400784B102851F6E21AC47090F8148E304C941D8CB13AD11343E17A971D8271949002C73",
		INITVAL_08 => "0x03A651162509CF915A0B102CD0F2460A2DC090C0170CB1148A0C0A9094A7048841F8FC10E31024C0",
		INITVAL_09 => "0x096180A60B042361BE291F413042311E80211C9A1DE6C1189E1F4D20B46B1A4C8178DC16AA81F043",
		INITVAL_0a => "0x07C671AC9D0C2E10504F0D28C152560428B0B47E150B714C8C1D6CA1C4C80A0D8120B90F05219C4F",
		INITVAL_0b => "0x0E8681D2BF164151568C1EC121E4AD004B81FCE10C2AF068D91D0F0124FA01E101BEBC1F8D31D858",
		INITVAL_0c => "0x02E4111C781AE7017A8C10423080A31288D02AB80945612A4109A2619E820D86C1642E0F43812689",
		INITVAL_0d => "0x068DB180521A0311721209EC11842602C0507E170FC510783F174181B4151CAF21426F104AF0F6AB",
		INITVAL_0e => "0x0C8301127010A161568519AD204AB815052092F00309E02ECD1F49C0E4300E270126761FA10104D1",
		INITVAL_0f => "0x0F8D814E020CADC1A09C0DA38030B60E07E0861401A230066D0A2AC1361C14A10080FE04A620745E",
		INITVAL_10 => "0x194AE0164A13E290E24F118B408C4D0485E1525416EE10300A1BC4D146AB0CA861EC3E00C9B0C097",
		INITVAL_11 => "0x09258080631F6491AC65156E01E094196DF0360B090A11C00E0E6350362B08A9E1F0AD17E471F885",
		INITVAL_12 => "0x0301506ECD120F2196A90C8390D690192BD0642C126EB0B0E21F00E194961B2521261A0D21414AB9",
		INITVAL_13 => "0x0BEE80208B17A101348E00CE7116ED0FC3806CED17EDE1644E1646C1D25C0A4300B88E128D810C42",
		INITVAL_14 => "0x024691D8601A02F1C29E0C41F1D2161E8411468216A17008BF17A0D0C84004683046E10FAA111843",
		INITVAL_15 => "0x1BE50116A6134ED0804D1C8EC1F21A114151B226090D71D2A519CC30B8841C2650203C1DE311B22F",
		INITVAL_16 => "0x1DE710B0A80D4E21F25B1B08A102A1020600DA83030160CE0215E4A1909519E2801A4E0B0BF0C860",
		INITVAL_17 => "0x10ADB08AFD046E016E23086A71E007134870BEB915E2B08C980C45815CE5156E41C8D40C6EA04E2F",
		INITVAL_18 => "0x0D6F8094120F485064D014E041189A10A58070900344F0D2A41E2D9018A31F4B80E20302A761AC74",
		INITVAL_19 => "0x0186A148761C4D41288318AF1086C3138541E4D2178F80F860042360C8C801A290644A072A71DE48",
		INITVAL_1a => "0x1D6531EAB2036CB1DAAF1AC2007A2B1503219696142591C015152E80C8FD17E0A146AE0EC501AE53",
		INITVAL_1b => "0x096B91145A0FA6802E6418E9A0863900240090A8030EB168B814E8B14A8B058B70089C0E09D1FAC2",
		INITVAL_1c => "0x1940F08C671A8EF1D2521848A078DB1384F0501D18C0C180D4192BA19AD014AA01928B1A41B15AEA",
		INITVAL_1d => "0x0E2121C2D4036E8194270A6530F4051E24F0B63D15ABF184FB01818170341B01E17E82130F907AB1",
		INITVAL_1e => "0x1040E0E0C00C2420E08B108C010892040141185E08EB0092870A6380B8A5138D71C289062541409A",
		INITVAL_1f => "0x0DE7619CC00F80D104261E6481D22005E210808B1B41012E4F07E820DE1D112BD14A8B1647A182CD",
		INITVAL_20 => "0x16A0703CED03C7E160ED01ABF1D0120D8620401A0388D04E010F8FA15CF60F0D10382109E0C0065E",
		INITVAL_21 => "0x052BC13E4805857170B6008CF0485C1365E060E20286B08E8F16A040D4831F0D416C6F18C2405AE0",
		INITVAL_22 => "0x0044315A46182FD07EB6136AB0180B10C541948E094350029F19CC81DA90074C8008F9162ED1DE82",
		INITVAL_23 => "0x0E476030AB174CE0CEBE092DB0C8060040A0E4FD040A40A06F1C47213EF30D6D012C321DAA818C27",
		INITVAL_24 => "0x194A40B6231242605E161E49D05031046C70E40B1C6870DE011863A0D6740C01E11231104D703A1F",
		INITVAL_25 => "0x0C8050206A0EA0B1F4A01CE1E1CEDE16414102FA186E7034BF0382B1A698158EF0BC1A1AEDE0683A",
		INITVAL_26 => "0x050700582518AE4164B2168B0050121F0C9080DC1A08E0562919CB61A202028751E21A18AD10025A",
		INITVAL_27 => "0x1E2A30AE5205E490861C08AF0138EC14C48140401F8D91F25A09E8C112D91E4B10D03C04E5A12C3D",
		INITVAL_28 => "0x19E180181C0F243014541D27D0161B0CAA009E46060A302AB81823D0C6780A8CE1DE981EC3A19C9D",
		INITVAL_29 => "0x0C441116720A6E80F2721B8E01D8950E0DC1CE141A0DF00E3F148EB0721B0906D108730484811806",
		INITVAL_2a => "0x1A04B1E6A00489705EAE070A0024241C6B61CED10B0CF196671465B114E90C8E8030321A8D917C62",
		INITVAL_2b => "0x1482F00EB808AD40701E0B05F0F2E10F83E1B023186D8126A60E4DC10C401CAF6052F91E2570460A",
		INITVAL_2c => "0x0583D13E18004FC162B418AFD012D61C687048F5142BD0BE390F4DE1C4171E840028B10D6DA196F0",
		INITVAL_2d => "0x1BCE71FA3F12CEA008B404EAD1FAB90D00C0E2EB0166D0D47C1705801C160788F148581F6280C67D",
		INITVAL_2e => "0x0B6BC1B49B0B20B08EBA180A91A6DE19CE20BE0C1608A048920E62F13E7A03CE302E86078AE1843C",
		INITVAL_2f => "0x0EC401BC7302A7A1267C1C87C15E2715A64138F619005140FC15E1405AA80746900E41090850FA37",
		INITVAL_30 => "0x0B0D70E84B0E47C10EA006EA3168B813E151FC0C0CA1714E151849B1802D112820BEA600636004D6",
		INITVAL_31 => "0x13C740F86712AAB18A3D02E310AE610CE42150520C4691147C1EACD15A83082AB0A6B80B8281E4F4",
		INITVAL_32 => "0x0E2BA01ECA10C28152CD04E5F03ECF0ECE415C7C1B02D180611FA3409CE11E4140423212E2E042F0",
		INITVAL_33 => "0x1BC451E2E30C8411E0E2190C11145F1900D142A1080760825309C061D25901E140C8AC1CED31BE94",
		INITVAL_34 => "0x080450B43D0DE460B0F40AE310462C064B803EC900CFB1B6A109EC61D2D91FCAF17CAE0A04A05C42",
		INITVAL_35 => "0x17EA0096E81606819A2410E7C05A52174C90E290060140EA1A0C2D4030311D0AD12EC3194B9064A7",
		INITVAL_36 => "0x1CADE0063C0E04D1C896086CB08EC0096901C6610E83A0DE8601CC81BE8E0F26C1C6050EA651F8DE",
		INITVAL_37 => "0x168BF02ABA1B8A3184E1194B21CE0A074F9064761C22300E7E0266006229064FE1C2241A4D21A678",
		INITVAL_38 => "0x0D2A7090DC1640D1AC5F1389C040A51B45A01E0B140A31C23C126A009A1F1641A1906C170AD14ED0",
		INITVAL_39 => "0x1FC6C026D708E170A42D16EB702AC50584D1305E14C14052FC0C65B19C971A87A1208A0BEA605003",
		INITVAL_3a => "0x17A7D074C1006EB020AD09069160AB114100A6371E0BC03E9714C261C8F808EEA134401EAE40E4F5",
		INITVAL_3b => "0x06AE2092B215A3C0507B14E32068C60528A0BEC8024231402E1704B16ABE09C70148460A8C701C9A",
		INITVAL_3c => "0x0C62507A350E8CF1205F0B24908C070C81A05ACF052960FA0115E7818C4F0180D10C0D006B501281",
		INITVAL_3d => "0x1C09613A2D0724E02E0D1B2071421D040B00A42018ABC17E650388B038ED020E50DA591CA1513E12",
		INITVAL_3e => "0x17CAD0B4611C6970607B1729405C15016691FC4219075128270E47611E50078CA1524A026C70DEDB",
		INITVAL_3f => "0x164D308A49116FB0A8131B6A3090411C61A1700A17CF0180E3038690A4D30EC790C0B909C9E1E6BA"
	)
	port map (
		DIA0 => '0', DIA1 => '0', DIA2 => '0', DIA3 => '0',
		DIA4 => '0', DIA5 => '0', DIA6 => '0', DIA7 => '0',
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => data_b(8), DOA1 => data_b(9),
		DOA2 => data_b(10), DOA3 => data_b(11),
		DOA4 => data_b(12), DOA5 => data_b(13),
		DOA6 => data_b(14), DOA7 => data_b(15),
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0', ADA2 => '0', 
		ADA3 => addr_b(2), ADA4 => addr_b(3),
		ADA5 => addr_b(4), ADA6 => addr_b(5),
		ADA7 => addr_b(6), ADA8 => addr_b(7),
		ADA9 => addr_b(8), ADA10 => addr_b(9),
		ADA11 => addr_b(10), ADA12 => addr_b(11),
		ADA13 => addr_b(12),
		CEA => '1', CLKA => clk_25m, WEA => '0',
		CSA0 => '0', CSA1 => '0', CSA2 => '0', RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => data_a(8), DOB1 => data_a(9),
		DOB2 => data_a(10), DOB3 => data_a(11),
		DOB4 => data_a(12), DOB5 => data_a(13),
		DOB6 => data_a(14), DOB7 => data_a(15),
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0', ADB2 => '0', 
		ADB3 => addr_a(2), ADB4 => addr_a(3),
		ADB5 => addr_a(4), ADB6 => addr_a(5),
		ADB7 => addr_a(6), ADB8 => addr_a(7),
		ADB9 => addr_a(8), ADB10 => addr_a(9),
		ADB11 => addr_a(10), ADB12 => addr_a(11),
		ADB13 => addr_a(12),
		CEB => '1', CLKB => clk_25m, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	ram_8_2: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B => "NORMAL", WRITEMODE_A => "NORMAL",
		GSR => "ENABLED", RESETMODE => "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A => "NOREG",
		DATA_WIDTH_B => 9, DATA_WIDTH_A => 9,
		INITVAL_00 => "0x1B413016D3112150823803EA91A88B0E6B00C6AE018611C42F0B2EA11C270E2120929E11ED807E06",
		INITVAL_01 => "0x0C297020FE0FC411A44F0DE4B01EE81EC3605A2005AD40DA2F1829C1E04817CD81246206C2D1CE37",
		INITVAL_02 => "0x002451DE1505060178CF0B276002F209ACF160E704E860B0F81F4E00F001078F8194700381E12A83",
		INITVAL_03 => "0x1FAF807C0E1F6A5138AC056210BCE400A9404AF51E4A313E8908C8F0722D1FCE91F0630406509E06",
		INITVAL_04 => "0x0D69A0DA3F0B6A61C84F06C290A882178E4102C813CB019C5215E20162EF196E41D0D40063A1BE25",
		INITVAL_05 => "0x070C30905C0EC8917A10140F01FAE51F02605A89028040D68B1FC0A0BCB7156D8126091E6581782B",
		INITVAL_06 => "0x1628A0E45A19224062980C44A006621E47B1A2D915A6105E620DA740566B1642B1926F0080E16826",
		INITVAL_07 => "0x0460F0CE2F0A2D90BEC2182D9026281E2BE0064A1806B012670E6FB0C675024BD11E5812EBE14A58",
		INITVAL_08 => "0x058FA05AEB05AD008CC70B69F004B006EFA0E6DB03C520F8D102ACF0D04517C9516401192CF19E67",
		INITVAL_09 => "0x0AEBD04CC2018870D4F61D2270965E04674078D813AD30D65A1C2390D2750186D03A7111EF41D4F5",
		INITVAL_0a => "0x19E1B186481F45A07A9A146FE0C8071A8F40EC14082AE1726D0E4F51E0BA046B907E50158FC1B298",
		INITVAL_0b => "0x1B2A50F06C09CFA01A5B164F01160E12A5E1A2B80189D1308F1FA1A08A5002CAF0C6D10C6E91369B",
		INITVAL_0c => "0x104A306E6A07843190960788F1BC460E42106CAC1F0C7056F21647011A1B042F00C85309A721B8B6",
		INITVAL_0d => "0x1A2EC1D63E18E7E0ECF6102F212E53078FC158050A0360D48C19E2711246112BC1C05119AB1048F9",
		INITVAL_0e => "0x13EDE0ECC6058FB1A2F2112B40E2651DA011B63409E470ACEA062761CA960A0BC11438194351D2B0",
		INITVAL_0f => "0x1A4EA172741E81A13EAB0821D0A6901B8AD1422B07E151F429064F10ECFD0C2EA0CEB9108CF1D078",
		INITVAL_10 => "0x1E2C709ABD0B0050CAA6074180E2820064A1F6100C4CF19A151F83809AE40F4DC112A112A260262D",
		INITVAL_11 => "0x1A47E0D2C202C8B106740D2A71AC230D2010A46D15AC007E240C4A91585C16435082F612A1505046",
		INITVAL_12 => "0x148FE1B4EB1F4C80046F012A70B47B0C4C7130700AE8C1264305C3D1A2C80D476158CF10EF013C40",
		INITVAL_13 => "0x0704A07A2405E4A078F30B88313E970585A002FA114030DE8F0E21B19E7A1EC940C6DB0A4CB0A6B0",
		INITVAL_14 => "0x0C6AB112231644317EF501E6C164BA156AD01AC909C8A03C5203479130DB0285701EA01D83013EE8",
		INITVAL_15 => "0x19C2314E1F018B40F4200A2A00804E0680E04C130BE1206AE11F0A701CB91A8271A4E2018A00846C",
		INITVAL_16 => "0x12668172F51B24F0B6C60E4760CAC814ED309E751A44808A610C88E03A04162560C88703E0A04E43",
		INITVAL_17 => "0x0F27E134961029C138761B29D0689A18E261048E168970E0261A8FC1B2100DA830E231002D1162DB",
		INITVAL_18 => "0x18AD91EAB61A2710EC370AC2E0524D0C4C315CC500E650046B074B602C8C06CA1040C6116A1048B6",
		INITVAL_19 => "0x16E891ECCB0EAA611C9E0FC6B0C28204A2B13CF31DA960CA7A19ADA13E3F1285403E780181509269",
		INITVAL_1a => "0x09EC01C28905EF20F84D194970400C0BCF50D25F1C8B6156F610C5A13EE01409E03AB91741A05004",
		INITVAL_1b => "0x0DA6D18EE1158C315A7501CDE0F47019A5A146C91CA950ECCA112650F6A61B2410A2A5184F81D815",
		INITVAL_1c => "0x016BE11ADB1461C05E4E01E5112A1707CB61A8EB1A67205E871BC7E0F4B2070951CE2409CEC01C98",
		INITVAL_1d => "0x0A46B00E7E040B40D08C1CEF01B03410C6915CE81E21A1D09C1B62E0E47E17CD8140370E88512472",
		INITVAL_1e => "0x07E5C0AC710EA561421507CBA1A4BF1BE5F1B203046A60F0260D04E11E0C11AB61067D0B406036D3",
		INITVAL_1f => "0x05A5C14EBA0306707C1703CB104059026460AC750F0A504A311DA7319A430589A092C10909605C92",
		INITVAL_20 => "0x1D02D050411F4420FCF904CDC17AC50121D072CD1D4470C82512CEC0E21D0ACA41B0BE024271F497",
		INITVAL_21 => "0x1D0A10A4D313EE21A2501F2BE0BE161EC1C03CFB1409F10CE312EAF0A021156861F45C0400710E97",
		INITVAL_22 => "0x196E7126511E481090C2084570E6E40FA010DAC21702915ECB162F30584F090231E40C0087404A71",
		INITVAL_23 => "0x0208C1EAE11A00A064FA06EE40E4490F69F1D6120EA061D2B401A0E0D69C02AAE07E01086D40B4B1",
		INITVAL_24 => "0x12603004EF1863F10272120C019EE519A8D17816158B51B2B403E180B8031828C148E80FCA0060DA",
		INITVAL_25 => "0x016B11D4781D4F5102C510A480368A0F05B0EAD90FA0307A6004CD6158650169C06E7E1D0FC12C86",
		INITVAL_26 => "0x0B89D0F2870569003AEC0E464128E41927313AB214C9C1C85C06AA01141C0BCB90C6650E22E0FA3F",
		INITVAL_27 => "0x1146D0D097116E20CE6D1E2CB00E1A1085903AD21B4601683614C161AEEF0B0E41F827168B701AC2",
		INITVAL_28 => "0x156BC1BC6706A1706CBA114E8094F6126C61B4D718C070D0F60C47214E320367B1B23701A4F1A0A8",
		INITVAL_29 => "0x0020A0D2100F497074D90367D0566305C28074070FC13168900B6CF0D82D1E23003649016FB162CF",
		INITVAL_2a => "0x08E2511C3D072821C29F12EB41B870094AC152CB052B91A0A30B27A1A2AF1B62C16AE8020B00E875",
		INITVAL_2b => "0x1EC5B0A67112EBF0B2D7024EC014741BC4004E5C1E043180811A2291F6210022B18A650782600AC1",
		INITVAL_2c => "0x030E210CF308CB10FAD910C240468A0F26312ECE170AF008761609C182CD10AD90A0070504B1FCE1",
		INITVAL_2d => "0x052C309248056B71D48D1B2831306A0949A0505C0BC9C1069014C711A48F11EE2036F90BC530026C",
		INITVAL_2e => "0x0D2E0120D8178EA026E80363C0FC2C1020416C721A2570AC741C8D80B69404ED700ABD03E781267A",
		INITVAL_2f => "0x072AD126481C89514E610B20B118E91181D1EC210747C08E85170A316EF413845172530FA3A1149A",
		INITVAL_30 => "0x1862E04C501BC2B056FD02A79114A40B8CB1A2F115EEC1DA4201A4013668048E30460C058C50F838",
		INITVAL_31 => "0x0E00B174BC1E4D8150C7168CD1C0C00627608A671F63402A13042711D85716E7C14065160B60B25A",
		INITVAL_32 => "0x07A7E1586D0E8B907C17162620D4A50A0D81B28604C6F126041566F1205719A6F178E1096B81B83E",
		INITVAL_33 => "0x072B8168C814EE3056340AE50162600BEBC180D70C49B14E68172D109020192BE07A0B0847C024E7",
		INITVAL_34 => "0x0B6FE072EC04858034E1040E81B27B11CEA178620388201C4701CD815074052060F27905CF3180B7",
		INITVAL_35 => "0x1B2DF134450F2BC02C3014C15162361B0FA1D6E318C3D062B706A7809CF21341418C2610A720CE3D",
		INITVAL_36 => "0x0263C0A2F6174200A07313A96106DE0422E0A28501C87134F317EF5174C917C101A8970D0A116434",
		INITVAL_37 => "0x152961580C0FC151E0DC12041172571D0C51E2D31F0601581D0BCC30A06F19A48180700923912CEC",
		INITVAL_38 => "0x1A86314E96118290586915E780728703E6C0ACF203874056F905C6C15C2310EDE12A2104EF611AFA",
		INITVAL_39 => "0x096091AEC612CA3170F6180180949800C6F16AA000E6A17ADA15271146C8064341DAC106CC80962E",
		INITVAL_3a => "0x1F4E41A8AF1E8941AEE71F2B71DA071283A0825E0C2861A6650F2B9160340B40306E6B0D47B162E4",
		INITVAL_3b => "0x1901D0FC010808A06A15080E50C4A708CD60469A10CED0CA8708C9E1D8CF030AD16EFA026851E260",
		INITVAL_3c => "0x11E9E050E20B28504A830E40302E6210676112530F04A1404E08C1B074B50EC72034AB0B49F04AE4",
		INITVAL_3d => "0x02E250689408AFA1B8C71CEA9196F81924A1EC3E0D67A084480E6250D0B11CE70072EB06EB8106B7",
		INITVAL_3e => "0x0BE841DEAD1B0DA0E4DE1CE871E80F03882124160C6C60C014092530B66901CDE08E3E04C1516240",
		INITVAL_3f => "0x09E7916C851820614E021086D1A6F61A8E81F4E51F82612CA8106DC0E2FC07202036EA10E7D15AC0"
	)
	port map (
		DIA0 => '0', DIA1 => '0', DIA2 => '0', DIA3 => '0',
		DIA4 => '0', DIA5 => '0', DIA6 => '0', DIA7 => '0',
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => data_b(16), DOA1 => data_b(17),
		DOA2 => data_b(18), DOA3 => data_b(19),
		DOA4 => data_b(20), DOA5 => data_b(21),
		DOA6 => data_b(22), DOA7 => data_b(23),
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0', ADA2 => '0', 
		ADA3 => addr_b(2), ADA4 => addr_b(3),
		ADA5 => addr_b(4), ADA6 => addr_b(5),
		ADA7 => addr_b(6), ADA8 => addr_b(7),
		ADA9 => addr_b(8), ADA10 => addr_b(9),
		ADA11 => addr_b(10), ADA12 => addr_b(11),
		ADA13 => addr_b(12),
		CEA => '1', CLKA => clk_25m, WEA => '0',
		CSA0 => '0', CSA1 => '0', CSA2 => '0', RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => data_a(16), DOB1 => data_a(17),
		DOB2 => data_a(18), DOB3 => data_a(19),
		DOB4 => data_a(20), DOB5 => data_a(21),
		DOB6 => data_a(22), DOB7 => data_a(23),
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0', ADB2 => '0', 
		ADB3 => addr_a(2), ADB4 => addr_a(3),
		ADB5 => addr_a(4), ADB6 => addr_a(5),
		ADB7 => addr_a(6), ADB8 => addr_a(7),
		ADB9 => addr_a(8), ADB10 => addr_a(9),
		ADB11 => addr_a(10), ADB12 => addr_a(11),
		ADB13 => addr_a(12),
		CEB => '1', CLKB => clk_25m, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	ram_8_3: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B => "NORMAL", WRITEMODE_A => "NORMAL",
		GSR => "ENABLED", RESETMODE => "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A => "NOREG",
		DATA_WIDTH_B => 9, DATA_WIDTH_A => 9,
		INITVAL_00 => "0x1C60C1E89608EE314E9C0560C1C0A1194650E48D13C3A08A931FC81182CD1B08607AA3196471527B",
		INITVAL_01 => "0x17A5E0B420186DB062DE09A5A0D6FB0749D1E6E40F829026160CAEB0862F1842F1AE49142460145C",
		INITVAL_02 => "0x18CBA186F21AC95052601968A15CC00641E18A810D01A084560BCB91743204AC3172D614E850905A",
		INITVAL_03 => "0x1023103AF90D40F0F43500A3C15895042DA1686A0BC94080A700EE414CF00A8DF1385909C81024DB",
		INITVAL_04 => "0x00AF6058961EC310B45B1924B1465F1D0810B661180241B438086F90DA521507D04E7B09E7E134B0",
		INITVAL_05 => "0x09ED8062F2182C213C5E1C61B1C6F21B4951F8CF1F05904E9E052960728A19032118E41A42F00CC5",
		INITVAL_06 => "0x0DEDB116EC146130B04200EDF034D01B01600EFC108D3086851060B0C84508A1010ACA1D2F302450",
		INITVAL_07 => "0x0802C0A8530DE8E1C639050CB0E0ED046291FC710BE500B6AD004621BEC90DE68126C916A541709A",
		INITVAL_08 => "0x0C04903C791F2A303E650E43817A7508C610CAAE084160ACCE184580A2E013A2E1B2620B4D611A39",
		INITVAL_09 => "0x1C446120F51CA5C1203C0A85E1A0741D0951AEB7056211244B06A0E06E210DE271F438038E90B2AE",
		INITVAL_0a => "0x034D8140FA09ABF13EED118A51BEA90602D120281ECC91A09F1A0E119A6F1E8A7184FC0D2EB0F46A",
		INITVAL_0b => "0x014931582900AB01C879102D41C89308CA9104F21AE3405A360425300E4115AC3140EA024420FA2F",
		INITVAL_0c => "0x0C68719AD30D25205E5F0A264172751B04E040E916C1B0CE0D130410C44E07EB9020F00C2151DEFC",
		INITVAL_0d => "0x0C4720AECF0620D0A050056361168C11AEA1DA2B0820A112D9030BC19C02194ED0E82006C58012E4",
		INITVAL_0e => "0x116CF1569212C8408C1E0CE170784F028CB0DE5915A3D1800F1C8B501272078620AECA016AC19EA7",
		INITVAL_0f => "0x0D6730B069124B018CE515EF414C5A1269B1BE681C26709CBC08E5615A600E637172AD1D6090AEC2",
		INITVAL_10 => "0x1BC830D27E194E3140D302EED07A9E0CE731C02B0808214664156F90E00D1803A07AD0156071EA8C",
		INITVAL_11 => "0x0DEC11A4591B4650348201E31046FE1504608C1216C750A4BD10A781BE171CEF01B4840D03212A1B",
		INITVAL_12 => "0x1D6BC1C0290D6930FA03174061805C0F6610FAB509C2518C1D1A2A71FCDA178401C0ED1566517825",
		INITVAL_13 => "0x182FB1841E012D30FA2D02E9D1942311246048BC1CA721A29B1BC5706406190FD150A701C2F04E6D",
		INITVAL_14 => "0x00A7C1E6541D20E14AA80B2820E85C0A0F609E6D0F4BE1A4980806C0F6210CEE418ACD120E507CA9",
		INITVAL_15 => "0x0464F0B85C0BC170363F0F09D0A40D1FAA41864F0C6401F4B702A05124DF11EB41F605162DC1FC10",
		INITVAL_16 => "0x01A5A1944E11683158F21D83D09457196F21129E1965F1465B0B09B17EEF0C0C9136310D4D101AD7",
		INITVAL_17 => "0x0788C0DE8C0CE5B14A8411E4B1C45E1703116C2F112601465F06E391907C11E790A62004E340A004",
		INITVAL_18 => "0x05262136D019024182A4008D30EC781827A182F307AB20B6890BCCA0A45E0A2EF08C950D8DC11EA9",
		INITVAL_19 => "0x04ADF1B21A1900F15A74164AC11AD717CE8008E91E2CB162D91FCC10646D0DE8F0D0BD15E4007A5A",
		INITVAL_1a => "0x002AF006760D8600261B0364B1286F072101E4280B0F202E401F8BC160390C2DF1C00C03A3F1922F",
		INITVAL_1b => "0x102C71620C160590809A04A8C1D0DC046930FCF61F4A0114651AC1408C1F0C6201D668036BC004FE",
		INITVAL_1c => "0x0EADA1E69403082008780B6E71F4A00A0A11F2F810E1B0AC26050D102C4F0D8F600A9E0022F196D4",
		INITVAL_1d => "0x00C8515A0B1DED703EE5138E9082691645208E471606402A500DED70281802EAB1D21C16CE411E0D",
		INITVAL_1e => "0x0D81F058B6046B81CA2F1E2F102648182861CE490125F1CA4503E1F12C3E1460A18E3E080FB1AE6C",
		INITVAL_1f => "0x092A30A09506C4B192CB1B47D08AFE0BCB70E4EA1864E1D66A12451062EA0EC0C06E2713AC80FA76",
		INITVAL_20 => "0x134C61F8B201A93158CB0E8161480B05AF318A6F1BEAE072B70505B060B8172FE1FC840A61D02C83",
		INITVAL_21 => "0x08EE0018711DA301F49715C580D28F09AB80EA840FA8D1241D04CD11E6E50282119A32172E912645",
		INITVAL_22 => "0x0D2180DEB21ACA415C0910C481C4D712627002D30D2480B6A61B4E11166203C1D0362D1BC39108E3",
		INITVAL_23 => "0x178D31488418E15080D911AA71B2AB13CD312A8C08CDB0E4820264D1B0E51E8F3114CF040BE1F004",
		INITVAL_24 => "0x01EEF182D00AC1406A0B0AC761C6780E0A101A2D02AAC150A61AC5E042D905A5F1B6421B6690F8C6",
		INITVAL_25 => "0x1AE2F0B8C9106AE19C371822F09A9B0D28F174BC02CC90C04117E7013CBF12C5A00230158A911ED9",
		INITVAL_26 => "0x026B401A6102EB51E8F10D2790AE301A60D0C69F0722B00AB01E4751C6E70E062058B71464818CC6",
		INITVAL_27 => "0x18AF9074C8082D01508A0166A0BCF507AEA08E6311C3701CF4002F51C8A406CFA13AD812A681F6F8",
		INITVAL_28 => "0x0D25E1E28A008601BE101BEB40FC0C0E831070311E2450F4241B096020E91D0981962E1649E16E6F",
		INITVAL_29 => "0x1B85E1B43C080B21D00B1D0C30BEC70363900ADE1346C1B42C0EC8D1E06F046711AC520CAEA0DAAB",
		INITVAL_2a => "0x1346F052410A0CB0B85C08A790E6611B017170F618C0212E980186817C8C0F013194D10E67E12ACB",
		INITVAL_2b => "0x00269058EA17C820DEC217C381A685114250781F0B49714CFC1088E058BD0E6590F0A00C4100ECDB",
		INITVAL_2c => "0x1C6F41742D16A2E1080E14E630BEC11184A1BC9B09A461D6A41A88A0160A0623A0D6420EA9F14A2B",
		INITVAL_2d => "0x10809164A900A0116A1F086940D60F0E2651BCA912E3A12ED31B23C1E8350B24B1CA6A1189409E32",
		INITVAL_2e => "0x05E2D0C62E1EC150D44905E650147915651148B519E63112BE1A4BE0D8B01B6020C8720DA490EA1D",
		INITVAL_2f => "0x1A8FB0945A064C80C0280E46A03C84026200703512E2E1CA1B02A8E0206500CBF1586A0C4171C20D",
		INITVAL_30 => "0x03E301A6A91706802A4609CE40DE6915086046530602B082E71C65A0DE9306EC70C0FB1BE9007271",
		INITVAL_31 => "0x1B6921C2D90864E12E6210CAF146A709A9503E1811AF80E8A619CE00264E0BC101EC9414CFD160BE",
		INITVAL_32 => "0x14CD417203172D410EE2018B806A9B094BF19E2B02EC10E47313C2814A4201C5201E850DACD1F09A",
		INITVAL_33 => "0x058921A4FD06AA51D8851C43A1F8A104C9E1AE0E1E2C516CC71EABA0A43F1D458112FE1B29E1D8A3",
		INITVAL_34 => "0x0D2980E0011623907EB01C2D419E5802E9D05A5306A6114E8E07473078B606015090030E61D02E50",
		INITVAL_35 => "0x05CBE00C1B14CF11E6F11A63619E790FCD3008A71FAEF09C64158121FA601E66B0A010136D010A10",
		INITVAL_36 => "0x0F481058A51B279146C2004FA02A1201C5F1842704A5C086DA05A291805A1B0AF052B4052F810A0A",
		INITVAL_37 => "0x01CC500E61024C703C021F65610AB90E2EB11CC00B6DC1A2381E4F20C8C300213146361F0061945B",
		INITVAL_38 => "0x0701402ABF0BC36130A00C0D31B89C068F8056410CE0600AAD1A81B1268D02C8C15CFD0B20108C69",
		INITVAL_39 => "0x01457104291A0561824B1426D17CBA1B2380ECB4162B711E3601EA411A2D11260058FD1823F1C29C",
		INITVAL_3a => "0x092BA0EC0614A7D08C300C4850E2CE0C6470CE48174FA14C2B11ACD02E6A026FC1BCFA018850ACA3",
		INITVAL_3b => "0x0CE831564F02E71082E21B6F10B29B0A0F401CB5186C016E590A4F203E980B4E112C531C0EB17853",
		INITVAL_3c => "0x0B44F1EC94006B60C869086F51A4391B4B50DE8908C3819CDB170561A016036E11F6EF08C2E196BA",
		INITVAL_3d => "0x18A031DE700D05B140E1068C31ACAC1F66F1164F050E500AB11D09705AF8094141F87C192C715805",
		INITVAL_3e => "0x092F9090B408EE40DA10150521A0CB1E44F1A0BF03AA81A4561A0411423F15ABF1A65918E320A471",
		INITVAL_3f => "0x1308A1F0FA0EA9D1C6CF0D4F814C3A012FC0D29F11A3115EDF1CAFA070160A06C0A4481460B12CF6"
	)
	port map (
		DIA0 => '0', DIA1 => '0', DIA2 => '0', DIA3 => '0',
		DIA4 => '0', DIA5 => '0', DIA6 => '0', DIA7 => '0',
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => data_b(24), DOA1 => data_b(25),
		DOA2 => data_b(26), DOA3 => data_b(27),
		DOA4 => data_b(28), DOA5 => data_b(29),
		DOA6 => data_b(30), DOA7 => data_b(31),
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0', ADA2 => '0', 
		ADA3 => addr_b(2), ADA4 => addr_b(3),
		ADA5 => addr_b(4), ADA6 => addr_b(5),
		ADA7 => addr_b(6), ADA8 => addr_b(7),
		ADA9 => addr_b(8), ADA10 => addr_b(9),
		ADA11 => addr_b(10), ADA12 => addr_b(11),
		ADA13 => addr_b(12),
		CEA => '1', CLKA => clk_25m, WEA => '0',
		CSA0 => '0', CSA1 => '0', CSA2 => '0', RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => data_a(24), DOB1 => data_a(25),
		DOB2 => data_a(26), DOB3 => data_a(27),
		DOB4 => data_a(28), DOB5 => data_a(29),
		DOB6 => data_a(30), DOB7 => data_a(31),
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0', ADB2 => '0', 
		ADB3 => addr_a(2), ADB4 => addr_a(3),
		ADB5 => addr_a(4), ADB6 => addr_a(5),
		ADB7 => addr_a(6), ADB8 => addr_a(7),
		ADB9 => addr_a(8), ADB10 => addr_a(9),
		ADB11 => addr_a(10), ADB12 => addr_a(11),
		ADB13 => addr_a(12),
		CEB => '1', CLKB => clk_25m, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

end x;
