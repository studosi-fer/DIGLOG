/* Verilog model created from schematic LV2.sch -- Nov 05, 2017 18:40 */

module LV2;




endmodule // LV2
